module mux8to1B32 (input logic C2,input logic C1, input logic C0, input logic [31:0] I3, 
	input logic[31:0] I2, input logic [31:0] I1, 
	input logic [31:0] I0, output logic [31:0] O);

	mux8to1B4 s1(C2,C1,C0,I7[3:0],I6[3:0],I5[3:0],I4[3:0],I3[3:0],I2[3:0],I1[3:0],I0[3:0],O[3:0]);
	mux8to1B4 s2(C2,C1,C0,I7[7:4],I6[7:4],I5[7:4],I4[7:4],I3[7:4],I2[7:4],I1[7:4],I0[7:4],O[7:4]);
	mux8to1B4 s3(C2,C1,C0,I7[11:8],I6[11:8],I5[11:8],I4[11:8],I3[11:8],I2[11:8],I1[11:8],I0[11:8],O[11:8]);
	mux8to1B4 s4(C2,C1,C0,I7[15:12],I6[15:12],I5[15:12],I4[15:12],I3[15:12],I2[15:12],I1[15:12],I0[15:12],O[15:12]);
	mux8to1B4 s5(C2,C1,C0,I7[19:16],I6[19:16],I5[19:16],I4[19:16],I3[19:16],I2[19:16],I1[19:16],I0[19:16],O[19:16]);
	mux8to1B4 s6(C2,C1,C0,I7[23:20],I6[23:20],I5[23:20],I4[23:20],I3[23:20],I2[23:20],I1[23:20],I0[23:20],O[23:20]);
	mux8to1B4 s7(C2,C1,C0,I7[27:24],I6[27:24],I5[27:24],I4[27:24],I3[27:24],I2[27:24],I1[27:24],I0[27:24],O[27:24]);
	mux8to1B4 s8(C2,C1,C0,I7[31:28],I6[31:28],I5[31:28],I4[31:28],I3[31:28],I2[31:28],I1[31:28],I0[31:28],O[31:28]);
	
endmodule
